** Profile: "SCHEMATIC1-D_Av_maxamp"  [ c:\cadence\my projects\lab_analogcad_exp4\lab_analogcad_exp4-PSpiceFiles\SCHEMATIC1\D_Av_maxamp.sim ] 

** Creating circuit file "D_Av_maxamp.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\sixsi\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1m 0 2u 
.STEP LIN PARAM Vamp1 100m 100m 100m 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
