** Profile: "SCHEMATIC1-freq_sweep"  [ d:\orcad projects\digi_elec_final9_v2\digi_elec_final9_v2-pspicefiles\schematic1\freq_sweep.sim ] 

** Creating circuit file "freq_sweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\sixsi\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 70m 60m 0.1u 
.STEP PARAM period LIST 1.05m 1.025m 1m 0.9m 0.8m 0.7m 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
