** Profile: "SCHEMATIC1-time_3stg"  [ D:\Orcad Projects\prep5_analog2_lab\prep5_analog2_lab-PSpiceFiles\SCHEMATIC1\time_3stg.sim ] 

** Creating circuit file "time_3stg.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\sixsi\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 3m 0 1u SKIPBP 
.STEP LIN PARAM pot_sweep 0 1.1 1 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
