** Profile: "SCHEMATIC1-prep_q3"  [ C:\Cadence\My projects\Lab_analogCAD_exp1\Lab_analogCAD_exp1-PSpiceFiles\SCHEMATIC1\prep_q3.sim ] 

** Creating circuit file "prep_q3.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\sixsi\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10m 0 10u 
.STEP LIN PARAM RVAL 50 4k 50 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
