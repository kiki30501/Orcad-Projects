** Profile: "SCHEMATIC1-HEHE"  [ D:\Orcad Projects\Diode_cap_calc\Diode_cap_calc-PSpiceFiles\SCHEMATIC1\HEHE.sim ] 

** Creating circuit file "HEHE.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../diode_cap_calc-pspicefiles/diode_cap_calc.lib" 
* From [PSPICE NETLIST] section of C:\Users\sixsi\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 0.5 0 1m 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
