** Profile: "SCHEMATIC1-circuit_3a_ampsweep"  [ c:\cadence\my projects\lab_analogcad_exp3\lab_analogcad_exp3-pspicefiles\schematic1\circuit_3a_ampsweep.sim ] 

** Creating circuit file "circuit_3a_ampsweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\sixsi\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1m 0 1u 
.STEP LIN PARAM Vamp 1.9 2.2 0.05 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
