** Profile: "SCHEMATIC4-2654"  [ d:\orcad projects\lab_dig_elec_5\lab_dig_elec_5-PSpiceFiles\SCHEMATIC4\2654.sim ] 

** Creating circuit file "2654.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\sixsi\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 2m 1m 1u SKIPBP 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC4.net" 


.END
