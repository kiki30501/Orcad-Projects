Library IEEE;