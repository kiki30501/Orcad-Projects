** Profile: "SCHEMATIC1-calc_1"  [ c:\cadence\my projects\lab_analogcad_exp1\lab_analogcad_exp1-PSpiceFiles\SCHEMATIC1\calc_1.sim ] 

** Creating circuit file "calc_1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../lab_analogcad_exp1-pspicefiles/lab_analogcad_exp1.lib" 
* From [PSPICE NETLIST] section of C:\Users\sixsi\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10m 0 100u 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
