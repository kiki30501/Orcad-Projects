** Profile: "SCHEMATIC1-circuit3a_DConly"  [ C:\Cadence\My projects\Lab_analogCAD_exp3\Lab_analogCAD_exp3-PSpiceFiles\SCHEMATIC1\circuit3a_DConly.sim ] 

** Creating circuit file "circuit3a_DConly.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\sixsi\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.OP
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
