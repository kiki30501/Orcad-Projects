** Profile: "SCHEMATIC1-dc_freq_sweep"  [ D:\Orcad Projects\digi_elec_final9\digi_elec_final9-PSpiceFiles\SCHEMATIC1\dc_freq_sweep.sim ] 

** Creating circuit file "dc_freq_sweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\sixsi\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 0.1 0 1u 
.STEP LIN PARAM {Period} 0.1 4.9 0.3 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
