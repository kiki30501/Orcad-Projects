** Profile: "SCHEMATIC1-q4a_without_body"  [ D:\Orcad Projects\hw5_dig_elec\hw5_digi_elec-PSpiceFiles\SCHEMATIC1\q4a_without_body.sim ] 

** Creating circuit file "q4a_without_body.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../hw5_digi_elec-pspicefiles/hw5_digi_elec.lib" 
* From [PSPICE NETLIST] section of C:\Users\sixsi\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_Vin 0 5 0.1m 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
