** Profile: "SCHEMATIC1-A_ID_VDS"  [ c:\cadence\my projects\lab_analogcad_exp4\lab_analogcad_exp4-PSpiceFiles\SCHEMATIC1\A_ID_VDS.sim ] 

** Creating circuit file "A_ID_VDS.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\sixsi\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V6 0 15 0.1 
+ LIN V_V1 0 5 0.5 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
